* SPICE3 file created from pass_or.ext - technology: scmos

.option scale=1u

M1000 B' inverter_0/in B' Gnd nfet w=8 l=2
+  ad=112 pd=72 as=0 ps=0
M1001 B' inverter_0/in B' B' pfet w=24 l=2
+  ad=304 pd=136 as=0 ps=0
M1002 VDD a_20_n12# a_12_n10# Gnd nfet w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1003 a_12_n10# B' a_2_n10# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=64 ps=32
C0 A Gnd 5.15fF **FLOATING
C1 B Gnd 5.38fF **FLOATING
C2 VDD Gnd 2.35fF
C3 a_20_n12# Gnd 3.81fF
C4 B' Gnd 22.14fF
C5 inverter_0/in Gnd 4.36fF
