magic
tech scmos
timestamp 1664280310
<< nwell >>
rect -9 -5 9 31
<< polysilicon >>
rect -1 21 1 23
rect -1 -14 1 -3
rect -1 -24 1 -22
<< ndiffusion >>
rect -7 -16 -1 -14
rect -7 -20 -6 -16
rect -2 -20 -1 -16
rect -7 -22 -1 -20
rect 1 -16 7 -14
rect 1 -20 2 -16
rect 6 -20 7 -16
rect 1 -22 7 -20
<< pdiffusion >>
rect -7 12 -1 21
rect -7 8 -6 12
rect -2 8 -1 12
rect -7 -3 -1 8
rect 1 12 7 21
rect 1 8 2 12
rect 6 8 7 12
rect 1 -3 7 8
<< metal1 >>
rect -15 34 17 39
rect -6 29 -2 34
rect -6 12 -2 25
rect 2 -16 6 8
rect -6 -25 -2 -20
rect -15 -26 17 -25
rect -15 -30 -6 -26
rect -2 -30 17 -26
<< ntransistor >>
rect -1 -22 1 -14
<< ptransistor >>
rect -1 -3 1 21
<< polycontact >>
rect -5 -11 -1 -7
<< ndcontact >>
rect -6 -20 -2 -16
rect 2 -20 6 -16
<< pdcontact >>
rect -6 8 -2 12
rect 2 8 6 12
<< psubstratepcontact >>
rect -6 -30 -2 -26
<< nsubstratencontact >>
rect -6 25 -2 29
<< labels >>
rlabel pdiffusion -5 -2 -5 -2 1 pdiffusion
rlabel ndcontact -4 -18 -4 -18 1 ndcontact
rlabel ndcontact 4 -18 4 -18 1 ndcontact
rlabel polycontact -3 -9 -3 -9 1 in
rlabel metal1 1 -28 1 -28 1 GND
rlabel metal1 4 -9 4 -9 1 out
rlabel nwell 2 25 2 25 1 nwell
rlabel nsubstratencontact -4 27 -4 27 1 nsubstratencontact
rlabel metal1 -1 36 -1 36 5 VDD
rlabel ptransistor 0 11 0 11 1 poly
rlabel pdcontact -4 10 -4 10 1 pdcontact
rlabel pdcontact 4 10 4 10 1 pdcontact
<< end >>
